`define TEST "hello"
    `define HELLO fun

"TEST __LINE__"

__LINE__ __FILE__ __DATE__ __TIME__

`define TEST2

`ifdef TEST2

`ifndef TEST4

TEST TEST TEST'test

"Hello there my name is TEST"

`else

tsktstk

`endif

TEST

`else

(TEST TEST: no TEST)

`endif

`ifndef TEST3

TEST TEST TEST_TEST HELLO

`endif

`define meow_1 "hello there my name is al"

meow_1
