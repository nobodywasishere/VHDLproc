`rand TEST1 B10

TEST1

`rand TEST2 D5

TEST2

`rand TEST3 H20

TEST3

`rand TEST4 A50

TEST4

`rand testing B1

testing
