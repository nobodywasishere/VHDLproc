`for 2

`for 4

`for 3

hello there

`endfor

`endfor

`endfor
