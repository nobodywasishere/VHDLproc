#define TEST2

#undef TEST2
