#for 10

hallo there

#endfor
