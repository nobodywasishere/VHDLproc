`if INCLUDE_FILE = 'true' then
`include '../tests/include-to.vhdl'
`else
`Warning "Not including thing"
`end if
