`include "include-to.vhdl"
