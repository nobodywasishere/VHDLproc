`define hello 4
`define there "people"

"hello there"
hello there
'hello there'
