`include '../tests/include-to.vhdl'
