`message This test was successful

`error this is an error message
