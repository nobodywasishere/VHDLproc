`include "include-to.vhdl"

this is a test
