`define TEST "hello"
`define HELLO fun

TEST


`define TEST2

`ifdef TEST2

`ifndef TEST4

TEST TEST TEST

`else

tsktstk

`endif

TEST

`else

TEST TEST no TEST

`endif

`ifndef TEST3

TEST TEST TEST HELLO

`endif
