#message "This test was successful"
