#include "include-to.vhdl"
