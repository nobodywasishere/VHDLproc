
`undef TEST3

TEST3

TEST2
