`if INCLUDE_FILE = "TRUE" then
`include '../tests/include-to.vhdl'
`else
`Warning "Not including thing"
`end if
