`if a = 'a' then
    `if b = 'b' then
        a = 'a' and b = 'b'
    `else
        a = 'a' and b /= 'b'
    `end
`end